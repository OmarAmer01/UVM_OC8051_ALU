// // ALU Assertions / Coverage

// module alu_ac (
//     alu_if _alu_if
// );
// property not_correct;
//   @(posedge _alu_if.clk) _alu_if.op_code |->
// endproperty
// endmodule
